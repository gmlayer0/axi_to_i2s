module axi2_to_i2s (
  input  wire        s_axi_ctrl_aclk   ,
  input  wire        s_axi_ctrl_aresetn,
  input  wire        s_axi_ctrl_awvalid,
  output wire        s_axi_ctrl_awready,
  input  wire [ 7:0] s_axi_ctrl_awaddr ,
  input  wire        s_axi_ctrl_arvalid,
  output wire        s_axi_ctrl_arready,
  input  wire [ 7:0] s_axi_ctrl_araddr ,
  input  wire        s_axi_ctrl_wvalid ,
  output wire        s_axi_ctrl_wready ,
  input  wire [31:0] s_axi_ctrl_wdata  ,
  output wire        s_axi_ctrl_bvalid ,
  input  wire        s_axi_ctrl_bready ,
  output wire [ 1:0] s_axi_ctrl_bresp  ,
  output wire        s_axi_ctrl_rvalid ,
  input  wire        s_axi_ctrl_rready ,
  output wire [31:0] s_axi_ctrl_rdata  ,
  output wire [ 1:0] s_axi_ctrl_rresp  ,
  output wire        irq               ,
  input  wire        aud_mclk          ,
  input  wire        aud_mrst          ,
  output wire        lrclk_out         ,
  output wire        sclk_out          ,
  output wire        sdata_0_out       ,
  input  wire        s_axis_aud_aclk   ,
  input  wire        s_axis_aud_aresetn,
  input  wire [31:0] s_axis_aud_tdata  ,
  input  wire [ 2:0] s_axis_aud_tid    ,
  input  wire        s_axis_aud_tvalid ,
  output wire        s_axis_aud_tready
);

endmodule